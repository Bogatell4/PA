
module Fetch(A,B,C);
input wire A,B;
output wire C;
endmodule