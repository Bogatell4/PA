
module Memory(

    );
endmodule
