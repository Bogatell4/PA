module fullsystem();
//wire input1, input2, result;
//Fetch Fetch32(input1,input2,result);
endmodule

//hello this is a test