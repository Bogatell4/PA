
module WriteBack(

    );
endmodule
