

module Decode (

/*inputs:


*/


);

endmodule