
//module for implementing the kyber algorithm

module Kyber(

    );
endmodule
