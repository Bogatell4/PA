
//this moduleis meant to include all the stages of the pipeline connected together


module fullsystem();
//wire input1, input2, result;
//Fetch Fetch32(input1,input2,result);
endmodule

