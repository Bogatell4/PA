
module Memory(
    input wire enable,
    input wire clk,
    input wire [4:0] dst,
    input wire [31:0] data_in,
    output reg [31:0] data_out
    );
    
    
    //reg []memory[]
    
    
endmodule
