
module Writeback(

    );
endmodule
